
// Ethernet_IP_TX.sv


